module Counter(MClock, Resetn, n);
	input MClock;
	input Resetn;
	output [3:0] n;
	
	


endmodule